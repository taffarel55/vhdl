
--EXEMPLO DE RAM


LIBRARY IEEE;
    USE IEEE.STD_LOGIC_1164.ALL;
    USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY RAM_TB IS 
-- empty
END ENTITY;

ARCHITECTURE BEV OF RAM_TB IS

SIGNAL DATAIN : STD_LOGIC_VECTOR(7 DOWNTO 0):="00000000";
SIGNAL ADDRESS : STD_LOGIC_VECTOR(7 DOWNTO 0):="00000000";
SIGNAL W_R : STD_LOGIC:='0';
SIGNAL DATAOUT : STD_LOGIC_VECTOR(7 DOWNTO 0);

-- DUT component
COMPONENT RAM IS
    PORT(DATAIN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
         ADDRESS : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
         W_R : IN STD_LOGIC;
         DATAOUT : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
         );
END COMPONENT;

BEGIN

  -- Connect DUT
  UUT: RAM PORT MAP(DATAIN, ADDRESS, W_R, DATAOUT);

  PROCESS
  BEGIN
    -- Write data into RAM
    WAIT FOR 100 ns;
    ADDRESS<="10000000";
    DATAIN<="01111111";
    WAIT FOR 100 ns;
    ADDRESS<="01000000";
    DATAIN<="10111111";
    WAIT FOR 100 ns;
    ADDRESS<="00100000";
    DATAIN<="11011111";
    WAIT FOR 100 ns;
    ADDRESS<="00010000";
    DATAIN<="11101111";
    WAIT FOR 110 ns;

    -- Read data from RAM
    W_R<='1';
    ADDRESS<="00000000";
    WAIT FOR 100 ns;
    ADDRESS<="10000000";
    WAIT FOR 100 ns;
    ADDRESS<="01000000";
    WAIT FOR 100 ns;
    ADDRESS<="00100000";
    WAIT FOR 100 ns;
    ADDRESS<="00010000";
    WAIT FOR 100 ns;
    
    ASSERT FALSE REPORT "Test done. Open EPWave to see signals." SEVERITY NOTE;
    WAIT;
  END PROCESS;

END BEV;
